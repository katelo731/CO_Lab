//Subject:     CO project 3 - Sign extend
//--------------------------------------------------------------------------------
//Version:     3.5
//--------------------------------------------------------------------------------
//Writer:      0513311 Lo Wen-Huei
//--------------------------------------------------------------------------------
//Date:        2018 / 5 / 21
//--------------------------------------------------------------------------------
//Description: extend sign bit of data_i to [31:16]data_o
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
);
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
wire    [16-1:0] data_i;
reg     [32-1:0] data_o;

//Sign extended
always @(*) 
begin
	data_o <= {{ 16{data_i[15]} }, {data_i[15:0]}};
end

endmodule      
     