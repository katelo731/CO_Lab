//Subject:     CO project 3 - Adder
//--------------------------------------------------------------------------------
//Version:     3.5
//--------------------------------------------------------------------------------
//Writer:      0513311 Lo Wen-Huei
//--------------------------------------------------------------------------------
//Date:        2018 / 5 / 21
//--------------------------------------------------------------------------------
//Description: design for get pc_shift4 / branch_addr
//--------------------------------------------------------------------------------

module Adder(
   src1_i,
	src2_i,
	sum_o
);
     
//I/O ports
input  [32-1:0]    src1_i;
input  [32-1:0]	 src2_i;
output [32-1:0]	 sum_o;

//Internal Signals
wire   [32-1:0]	 sum_o;
//Parameter
    
//Main function
assign sum_o = src1_i + src2_i;

endmodule





                    
                    